/*  This file is part of JT6295.
    JT6295 program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    JT6295 program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with JT6295.  If not, see <http://www.gnu.org/licenses/>.

    Author: Jose Tejada Gomez. Twitter: @topapate
    Version: 1.0
    Date: 6-1-2020 */

// SS low  = divides by 164 (25.6 and 6.5kHz)
// SS high = divides by 132 (32   and 8  kHz)

module jt6295_timing(
    input       clk,
    input       cen,
    input       ss,
    output reg  cen_sr, // Sample rate
    output reg  cen_sr4 // 4x sample rate
);

reg  [2:0] base=2'd0;
reg  [5:0] cnt =8'd0;
wire [2:0] lim = ss ? 3'h3 : 3'h4;


always @(posedge clk) begin
    cen_sr4 <= 1'd0;
    cen_sr  <= 1'd0;
    if( cen ) begin
        base    <= (base==lim) ? 3'd0 : 3'd1;
        if(base==3'd0) cnt <= (cnt==6'd32) ? 6'd0 : cnt+6'd1;

        cen_sr4 <= ~base[2];
        cen_sr  <= {cnt,base} == 9'd0;
    end
end

endmodule
